-- Copyright (c) 2007-2020 Vitaly Chipounov
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

--------------------------------------------------
--UART Receiver
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.uart_lib.all;
use work.functions.all;

--To use the receiver, the clock speed parameter
--must be set to the frequency generated by the PLL.
--This generic parameter is used by the receiver to
--configure the internal counters to match the
--specified baud rate.
--This UART uses even parity.
entity uart_recv is
  generic (
    clock_speed : natural := 33000000;
    baud_rate : natural := 115200
  );
  port (
    clk : in std_logic;
    reset : in std_logic;
    --Receive connector on the board
    rx : in std_logic;
    --Asserted when a byte is received
    ready : out std_logic;
    --The received data
    data : out unsigned(7 downto 0);
    --Asserted when the parity of the received
    --byte is right.
    parity_ok : out std_logic
  );
end uart_recv;

architecture a1 of uart_recv is
  constant cc_size : natural := log2(clock_speed/baud_rate);
  signal rx_data_en : std_logic;
  signal sc_iseleven : std_logic;
  signal cc_incr : std_logic;
  signal cc_reset : std_logic;
  signal cc_max : unsigned(cc_size - 1 downto 0);
  signal cc_half : unsigned(cc_size - 1 downto 0);
begin
  dp : uart_recv_dp
  generic map(cc_size => cc_size)
  port map(
    clk => clk, reset => reset, rx => rx, data => data,
    rx_data_en => rx_data_en, sc_iseleven => sc_iseleven,
    cc_incr => cc_incr, cc_reset => cc_reset,
    cc_max => cc_max, cc_half => cc_half,
    parity_ok => parity_ok);

  sm : uart_recv_sm
  generic map(
    clock_speed => clock_speed, baud_rate => baud_rate,
    cc_size => cc_size)
  port map(
    clk => clk, reset => reset, rx => rx,
    ready => ready,
    rx_data_en => rx_data_en, sc_iseleven => sc_iseleven,
    cc_incr => cc_incr, cc_reset => cc_reset,
    cc_max => cc_max, cc_half => cc_half);

end a1;